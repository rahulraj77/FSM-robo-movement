localparam  IDLE      = 3'd0,
            FORWARD   = 3'd1,
            BACKWARD  = 3'd2,
            LEFT      = 3'd3,
            RIGHT     = 3'd4,
            STOP      = 3'd5,
            ERROR     = 3'd6,
            RECOVER   = 3'd7;
